//`timescale 1ns / 1ps
`include "ControlSignalDefine.v"
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/08/27 17:01:10
// Design Name: 
// Module Name: MemDataExtension
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module MemDataExtension(
    input [31:0] ReadMemData,
    input [3:0] ReadMemExtSignal,
    output reg[31:0] MemDataExt
    );
    
    always @(*) begin
      case (ReadMemExtSignal)
        `U_DWORD: MemDataExt = ReadMemData;
        `U_WORD_LOW: MemDataExt = {16'b0,ReadMemData[15:0]};
        `U_WORD_HIGH: MemDataExt = {16'b0,ReadMemData[31:16]};
        `U_BYTE_LOWEST: MemDataExt = {24'b0,ReadMemData[7:0]};
        `U_BYTE_LOW: MemDataExt = {24'b0,ReadMemData[15:8]};
        `U_BYTE_HIGH: MemDataExt = {24'b0,ReadMemData[23:16]};
        `U_BYTE_HIGHEST: MemDataExt = {24'b0,ReadMemData[31:24]};
        `S_WORD_LOW: MemDataExt = {{16{ReadMemData[15]}},ReadMemData[15:0]};
        `S_WORD_HIGH: MemDataExt = {{16{ReadMemData[31]}},ReadMemData[31:16]};
        `S_BYTE_LOWEST: MemDataExt = {{24{ReadMemData[7]}},ReadMemData[7:0]};
        `S_BYTE_LOW: MemDataExt = {{24{ReadMemData[15]}},ReadMemData[15:8]};
        `S_BYTE_HIGH: MemDataExt = {{24{ReadMemData[23]}},ReadMemData[23:16]};
        `S_BYTE_HIGHEST: MemDataExt = {{24{ReadMemData[31]}},ReadMemData[31:24]};
        default: ;
      endcase  
    end
    
endmodule
